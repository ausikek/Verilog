// 8-BIT REGISTER

`timescale 1ns/1ps
`include "combinational.v"

module reg8a (
        
    output wire [7:0] Reg_Out,
    input wire clk, res, EN,
    input wire [7:0] Reg_In
    
    );

    wire [7:0] nQ;
    wire [7:0] Mux_Out;

    MUX2_1 mux0 (Mux_Out, EN, Reg_Out, Reg_In);

    dflipflop dff0 (Reg_Out[0], nQ[1], clk, res, 1'b1, Mux_Out[0]);
    dflipflop dff1 (Reg_Out[1], nQ[0], clk, res, 1'b1, Mux_Out[1]);
    dflipflop dff2 (Reg_Out[2], nQ[3], clk, res, 1'b1, Mux_Out[2]);
    dflipflop dff3 (Reg_Out[3], nQ[2], clk, res, 1'b1, Mux_Out[3]);
    dflipflop dff4 (Reg_Out[4], nQ[5], clk, res, 1'b1, Mux_Out[4]);
    dflipflop dff5 (Reg_Out[5], nQ[4], clk, res, 1'b1, Mux_Out[5]);
    dflipflop dff6 (Reg_Out[6], nQ[7], clk, res, 1'b1, Mux_Out[6]);
    dflipflop dff7 (Reg_Out[7], nQ[6], clk, res, 1'b1, Mux_Out[7]);

endmodule